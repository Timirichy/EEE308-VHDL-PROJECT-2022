LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY STP_WTCH IS
PORT ( CLK50MHZ : IN  STD_LOGIC;
		 KEY      : IN  STD_LOGIC_VECTOR(1 DOWNTO 0);
		 SW       : IN  STD_LOGIC_VECTOR(9 DOWNTO 0);
		 LEDR     : OUT STD_LOGIC_VECTOR(9 DOWNTO 0);
		 HEX0     : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
		 HEX1     : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
		 HEX2     : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
		 HEX3     : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
		 HEX4     : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
		 HEX5     : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
		 );
END ENTITY STP_WTCH;


ARCHITECTURE behaviour OF STP_WTCH IS
SIGNAL CLK_play         : STD_LOGIC;
SIGNAL CLK_dis          : STD_LOGIC;
SIGNAL SEC_FLIP         : STD_LOGIC:='1';
SIGNAL MIC_SEC_FLIP     : STD_LOGIC:='1';
SIGNAL RSEST, STRT, STP : STD_LOGIC;
SIGNAL K                : STD_LOGIC := '0';
SIGNAL L                : STD_LOGIC := '1';
SIGNAL M                : STD_LOGIC_VECTOR(3 DOWNTO 0) := "0000";
SIGNAL N                : STD_LOGIC;

BEGIN

STRT             <=          KEY(0);
STP              <=          KEY(1);
RSEST            <=           SW(9);


DISP_CLK_3: WORK.Pl_CLK  PORT MAP(clk_3 => CLK50MHZ,
											T2     => CLK_play);
DISP_CLK_4: WORK.Dis_CLK PORT MAP(clk_4 => CLK50MHZ,
											T3     => CLK_dis);

PROCESS(CLK_play, CLK_dis, N, M, RSEST, MIC_SEC_FLIP, SEC_FLIP, STRT, STP, K, L)
VARIABLE P1, P2, P3 : INTEGER := 0;
BEGIN

	IF RISING_EDGE(CLK_dis) THEN
		IF M = "1011" THEN
			M <= "1011";
			N <= '1';
		ELSIF M /= "1011" THEN
			M <= M + "0001";
			N <= '0';
		END IF;
	END IF;
	
	
	
	IF N <= '0' THEN
		IF M <= "0000" THEN
			HEX0 <= STD_LOGIC_VECTOR'("10000110");
			HEX1 <= STD_LOGIC_VECTOR'("11111111");
			HEX2 <= STD_LOGIC_VECTOR'("11111111");
			HEX3 <= STD_LOGIC_VECTOR'("11111111");
			HEX4 <= STD_LOGIC_VECTOR'("11111111");
			HEX5 <= STD_LOGIC_VECTOR'("11111111");
		ELSIF M <= "0001" THEN
			HEX0 <= STD_LOGIC_VECTOR'("10000110");
			HEX1 <= STD_LOGIC_VECTOR'("10000110");
			HEX2 <= STD_LOGIC_VECTOR'("11111111");
			HEX3 <= STD_LOGIC_VECTOR'("11111111");
			HEX4 <= STD_LOGIC_VECTOR'("11111111");
			HEX5 <= STD_LOGIC_VECTOR'("11111111");
		ELSIF M <= "0010" THEN
			HEX0 <= STD_LOGIC_VECTOR'("10000110");
			HEX1 <= STD_LOGIC_VECTOR'("10000110");
			HEX2 <= STD_LOGIC_VECTOR'("10000110");
			HEX3 <= STD_LOGIC_VECTOR'("11111111");
			HEX4 <= STD_LOGIC_VECTOR'("11111111");
			HEX5 <= STD_LOGIC_VECTOR'("11111111");
		ELSIF M <= "0011" THEN
			HEX0 <= STD_LOGIC_VECTOR'("10110000");
			HEX1 <= STD_LOGIC_VECTOR'("10000110");
			HEX2 <= STD_LOGIC_VECTOR'("10000110");
			HEX3 <= STD_LOGIC_VECTOR'("10000110");
			HEX4 <= STD_LOGIC_VECTOR'("11111111");
			HEX5 <= STD_LOGIC_VECTOR'("11111111");
		ELSIF M <= "0100" THEN
			HEX0 <= STD_LOGIC_VECTOR'("11000000");
			HEX1 <= STD_LOGIC_VECTOR'("10110000");
			HEX2 <= STD_LOGIC_VECTOR'("10000110");
			HEX3 <= STD_LOGIC_VECTOR'("10000110");
			HEX4 <= STD_LOGIC_VECTOR'("10000110");
			HEX5 <= STD_LOGIC_VECTOR'("11111111");
		ELSIF M <= "0101" THEN
			HEX0 <= STD_LOGIC_VECTOR'("10000000");
			HEX1 <= STD_LOGIC_VECTOR'("11000000");
			HEX2 <= STD_LOGIC_VECTOR'("10110000");
			HEX3 <= STD_LOGIC_VECTOR'("10000110");
			HEX4 <= STD_LOGIC_VECTOR'("10000110");
			HEX5 <= STD_LOGIC_VECTOR'("10000110");
		ELSIF M <= "0110" THEN
			HEX0 <= STD_LOGIC_VECTOR'("11111111");
			HEX1 <= STD_LOGIC_VECTOR'("10000000");
			HEX2 <= STD_LOGIC_VECTOR'("11000000");
			HEX3 <= STD_LOGIC_VECTOR'("10110000");
			HEX4 <= STD_LOGIC_VECTOR'("10000110");
			HEX5 <= STD_LOGIC_VECTOR'("10000110");
		ELSIF M <= "0111" THEN
			HEX0 <= STD_LOGIC_VECTOR'("11111111");
			HEX1 <= STD_LOGIC_VECTOR'("11111111");
			HEX2 <= STD_LOGIC_VECTOR'("10000000");
			HEX3 <= STD_LOGIC_VECTOR'("11000000");
			HEX4 <= STD_LOGIC_VECTOR'("10110000");
			HEX5 <= STD_LOGIC_VECTOR'("10000110");
		ELSIF M <= "1000" THEN
			HEX0 <= STD_LOGIC_VECTOR'("11111111");
			HEX1 <= STD_LOGIC_VECTOR'("11111111");
			HEX2 <= STD_LOGIC_VECTOR'("11111111");
			HEX3 <= STD_LOGIC_VECTOR'("10000000");
			HEX4 <= STD_LOGIC_VECTOR'("11000000");
			HEX5 <= STD_LOGIC_VECTOR'("10110000");
		ELSIF M <= "1001" THEN
			HEX0 <= STD_LOGIC_VECTOR'("11111111");
			HEX1 <= STD_LOGIC_VECTOR'("11111111");
			HEX2 <= STD_LOGIC_VECTOR'("11111111");
			HEX3 <= STD_LOGIC_VECTOR'("11111111");
			HEX4 <= STD_LOGIC_VECTOR'("10000000");
			HEX5 <= STD_LOGIC_VECTOR'("11000000");
		ELSIF M <= "1010" THEN
			HEX0 <= STD_LOGIC_VECTOR'("11111111");
			HEX1 <= STD_LOGIC_VECTOR'("11111111");
			HEX2 <= STD_LOGIC_VECTOR'("11111111");
			HEX3 <= STD_LOGIC_VECTOR'("11111111");
			HEX4 <= STD_LOGIC_VECTOR'("11111111");
			HEX5 <= STD_LOGIC_VECTOR'("10000000");
		ELSE
			HEX0 <= STD_LOGIC_VECTOR'("11111111");
			HEX1 <= STD_LOGIC_VECTOR'("11111111");
			HEX2 <= STD_LOGIC_VECTOR'("11111111");
			HEX3 <= STD_LOGIC_VECTOR'("11111111");
			HEX4 <= STD_LOGIC_VECTOR'("11111111");
			HEX5 <= STD_LOGIC_VECTOR'("11111111");
		END IF;
	ELSE
		
		IF STRT = '0' AND STP = '1' THEN
			K <= '1';
			L <= '0';
		END IF;
		
		IF STP = '0' AND STRT = '1' THEN
			L <= '1';
			K <= '0';
		END IF;
		
		IF RISING_EDGE(CLK_play) THEN
					
			IF K <= '1' AND L <= '0' THEN
				IF RSEST = '1' THEN
					P1 := P1 + 1;
				ELSE
					P1 := 0;
				END IF;
			ELSIF K <= '0' AND L <= '1' THEN
				IF RSEST = '1' THEN
					P1 := P1;
				ELSE
					P1 := 0;
				END IF;
			END IF;
					
			IF (P1 = 100) THEN
				MIC_SEC_FLIP <= '0';
				P1 :=   0;
			ELSE
				MIC_SEC_FLIP <= '1';
				P1 :=   P1;
			END IF;
			
			IF P1 = 0 THEN
				HEX0 <= STD_LOGIC_VECTOR'("01000000");
				HEX1 <= STD_LOGIC_VECTOR'("11000000");
			ELSIF P1 = 1 THEN
				HEX0 <= STD_LOGIC_VECTOR'("01111001");
				HEX1 <= STD_LOGIC_VECTOR'("11000000");
			ELSIF P1 = 2 THEN
				HEX0 <= STD_LOGIC_VECTOR'("00100100");
				HEX1 <= STD_LOGIC_VECTOR'("11000000");
			ELSIF P1 = 3 THEN
				HEX0 <= STD_LOGIC_VECTOR'("00110000");
				HEX1 <= STD_LOGIC_VECTOR'("11000000");
			ELSIF P1 = 4 THEN
				HEX0 <= STD_LOGIC_VECTOR'("00011001");
				HEX1 <= STD_LOGIC_VECTOR'("11000000");
			ELSIF P1 = 5 THEN
				HEX0 <= STD_LOGIC_VECTOR'("00010010");
				HEX1 <= STD_LOGIC_VECTOR'("11000000");
			ELSIF P1 = 6 THEN
				HEX0 <= STD_LOGIC_VECTOR'("00000010");
				HEX1 <= STD_LOGIC_VECTOR'("11000000");
			ELSIF P1 = 7 THEN
				HEX0 <= STD_LOGIC_VECTOR'("01111000");
				HEX1 <= STD_LOGIC_VECTOR'("11000000");
			ELSIF P1 = 8 THEN
				HEX0 <= STD_LOGIC_VECTOR'("00000000");
				HEX1 <= STD_LOGIC_VECTOR'("11000000");
			ELSIF P1 = 9 THEN
				HEX0 <= STD_LOGIC_VECTOR'("00011000");
				HEX1 <= STD_LOGIC_VECTOR'("11000000");
			ELSIF P1 = 10 THEN
				HEX0 <= STD_LOGIC_VECTOR'("01000000");
				HEX1 <= STD_LOGIC_VECTOR'("11111001");
			ELSIF P1 = 11 THEN
				HEX0 <= STD_LOGIC_VECTOR'("01111001");
				HEX1 <= STD_LOGIC_VECTOR'("11111001");
			ELSIF P1 = 12 THEN
				HEX0 <= STD_LOGIC_VECTOR'("00100100");
				HEX1 <= STD_LOGIC_VECTOR'("11111001");
			ELSIF P1 = 13 THEN
				HEX0 <= STD_LOGIC_VECTOR'("00110000");
				HEX1 <= STD_LOGIC_VECTOR'("11111001");
			ELSIF P1 = 14 THEN
				HEX0 <= STD_LOGIC_VECTOR'("00011001");
				HEX1 <= STD_LOGIC_VECTOR'("11111001");
			ELSIF P1 = 15 THEN
				HEX0 <= STD_LOGIC_VECTOR'("00010010");
				HEX1 <= STD_LOGIC_VECTOR'("11111001");
			ELSIF P1 = 16 THEN
				HEX0 <= STD_LOGIC_VECTOR'("00000010");
				HEX1 <= STD_LOGIC_VECTOR'("11111001");
			ELSIF P1 = 17 THEN
				HEX0 <= STD_LOGIC_VECTOR'("01111000");
				HEX1 <= STD_LOGIC_VECTOR'("11111001");
			ELSIF P1 = 18 THEN
				HEX0 <= STD_LOGIC_VECTOR'("00000000");
				HEX1 <= STD_LOGIC_VECTOR'("11111001");
			ELSIF P1 = 19 THEN
				HEX0 <= STD_LOGIC_VECTOR'("00011000");
				HEX1 <= STD_LOGIC_VECTOR'("11111001");
			ELSIF P1 = 20 THEN
				HEX0 <= STD_LOGIC_VECTOR'("01000000");
				HEX1 <= STD_LOGIC_VECTOR'("10100100");
			ELSIF P1 = 21 THEN
				HEX0 <= STD_LOGIC_VECTOR'("01111001");
				HEX1 <= STD_LOGIC_VECTOR'("10100100");
			ELSIF P1 = 22 THEN
				HEX0 <= STD_LOGIC_VECTOR'("00100100");
				HEX1 <= STD_LOGIC_VECTOR'("10100100");
			ELSIF P1 = 23 THEN
				HEX0 <= STD_LOGIC_VECTOR'("00110000");
				HEX1 <= STD_LOGIC_VECTOR'("10100100");
			ELSIF P1 = 24 THEN
				HEX0 <= STD_LOGIC_VECTOR'("00011001");
				HEX1 <= STD_LOGIC_VECTOR'("10100100");
			ELSIF P1 = 25 THEN
				HEX0 <= STD_LOGIC_VECTOR'("00010010");
				HEX1 <= STD_LOGIC_VECTOR'("10100100");
			ELSIF P1 = 26 THEN
				HEX0 <= STD_LOGIC_VECTOR'("00000010");
				HEX1 <= STD_LOGIC_VECTOR'("10100100");
			ELSIF P1 = 27 THEN
				HEX0 <= STD_LOGIC_VECTOR'("01111000");
				HEX1 <= STD_LOGIC_VECTOR'("10100100");
			ELSIF P1 = 28 THEN
				HEX0 <= STD_LOGIC_VECTOR'("00000000");
				HEX1 <= STD_LOGIC_VECTOR'("10100100");
			ELSIF P1 = 29 THEN
				HEX0 <= STD_LOGIC_VECTOR'("00011000");
				HEX1 <= STD_LOGIC_VECTOR'("10100100");
			ELSIF P1 = 30 THEN
				HEX0 <= STD_LOGIC_VECTOR'("01000000");
				HEX1 <= STD_LOGIC_VECTOR'("10110000");
			ELSIF P1 = 31 THEN
				HEX0 <= STD_LOGIC_VECTOR'("01111001");
				HEX1 <= STD_LOGIC_VECTOR'("10110000");
			ELSIF P1 = 32 THEN
				HEX0 <= STD_LOGIC_VECTOR'("00100100");
				HEX1 <= STD_LOGIC_VECTOR'("10110000");
			ELSIF P1 = 33 THEN
				HEX0 <= STD_LOGIC_VECTOR'("00110000");
				HEX1 <= STD_LOGIC_VECTOR'("10110000");
			ELSIF P1 = 34 THEN
				HEX0 <= STD_LOGIC_VECTOR'("00011001");
				HEX1 <= STD_LOGIC_VECTOR'("10110000");
			ELSIF P1 = 35 THEN
				HEX0 <= STD_LOGIC_VECTOR'("00010010");
				HEX1 <= STD_LOGIC_VECTOR'("10110000");
			ELSIF P1 = 36 THEN
				HEX0 <= STD_LOGIC_VECTOR'("00000010");
				HEX1 <= STD_LOGIC_VECTOR'("10110000");
			ELSIF P1 = 37 THEN
				HEX0 <= STD_LOGIC_VECTOR'("01111000");
				HEX1 <= STD_LOGIC_VECTOR'("10110000");
			ELSIF P1 = 38 THEN
				HEX0 <= STD_LOGIC_VECTOR'("00000000");
				HEX1 <= STD_LOGIC_VECTOR'("10110000");
			ELSIF P1 = 39 THEN
				HEX0 <= STD_LOGIC_VECTOR'("00011000");
				HEX1 <= STD_LOGIC_VECTOR'("10110000");
			ELSIF P1 = 40 THEN
				HEX0 <= STD_LOGIC_VECTOR'("01000000");
				HEX1 <= STD_LOGIC_VECTOR'("10011001");
			ELSIF P1 = 41 THEN
				HEX0 <= STD_LOGIC_VECTOR'("01111001");
				HEX1 <= STD_LOGIC_VECTOR'("10011001");
			ELSIF P1 = 42 THEN
				HEX0 <= STD_LOGIC_VECTOR'("00100100");
				HEX1 <= STD_LOGIC_VECTOR'("10011001");
			ELSIF P1 = 43 THEN
				HEX0 <= STD_LOGIC_VECTOR'("00110000");
				HEX1 <= STD_LOGIC_VECTOR'("10011001");
			ELSIF P1 = 44 THEN
				HEX0 <= STD_LOGIC_VECTOR'("00011001");
				HEX1 <= STD_LOGIC_VECTOR'("10011001");
			ELSIF P1 = 45 THEN
				HEX0 <= STD_LOGIC_VECTOR'("00010010");
				HEX1 <= STD_LOGIC_VECTOR'("10011001");
			ELSIF P1 = 46 THEN
				HEX0 <= STD_LOGIC_VECTOR'("00000010");
				HEX1 <= STD_LOGIC_VECTOR'("10011001");
			ELSIF P1 = 47 THEN
				HEX0 <= STD_LOGIC_VECTOR'("01111000");
				HEX1 <= STD_LOGIC_VECTOR'("10011001");
			ELSIF P1 = 48 THEN
				HEX0 <= STD_LOGIC_VECTOR'("00000000");
				HEX1 <= STD_LOGIC_VECTOR'("10011001");
			ELSIF P1 = 49 THEN
				HEX0 <= STD_LOGIC_VECTOR'("00011000");
				HEX1 <= STD_LOGIC_VECTOR'("10011001");
			ELSIF P1 = 50 THEN
				HEX0 <= STD_LOGIC_VECTOR'("01000000");
				HEX1 <= STD_LOGIC_VECTOR'("10010010");
			ELSIF P1 = 51 THEN
				HEX0 <= STD_LOGIC_VECTOR'("01111001");
				HEX1 <= STD_LOGIC_VECTOR'("10010010");
			ELSIF P1 = 52 THEN
				HEX0 <= STD_LOGIC_VECTOR'("00100100");
				HEX1 <= STD_LOGIC_VECTOR'("10010010");
			ELSIF P1 = 53 THEN
				HEX0 <= STD_LOGIC_VECTOR'("00110000");
				HEX1 <= STD_LOGIC_VECTOR'("10010010");
			ELSIF P1 = 54 THEN
				HEX0 <= STD_LOGIC_VECTOR'("00011001");
				HEX1 <= STD_LOGIC_VECTOR'("10010010");
			ELSIF P1 = 55 THEN
				HEX0 <= STD_LOGIC_VECTOR'("00010010");
				HEX1 <= STD_LOGIC_VECTOR'("10010010");
			ELSIF P1 = 56 THEN
				HEX0 <= STD_LOGIC_VECTOR'("00000010");
				HEX1 <= STD_LOGIC_VECTOR'("10010010");
			ELSIF P1 = 57 THEN
				HEX0 <= STD_LOGIC_VECTOR'("01111000");
				HEX1 <= STD_LOGIC_VECTOR'("10010010");
			ELSIF P1 = 58 THEN
				HEX0 <= STD_LOGIC_VECTOR'("00000000");
				HEX1 <= STD_LOGIC_VECTOR'("10010010");
			ELSIF P1 = 59 THEN
				HEX0 <= STD_LOGIC_VECTOR'("00011000");
				HEX1 <= STD_LOGIC_VECTOR'("10010010");
			ELSIF P1 = 60 THEN
				HEX0 <= STD_LOGIC_VECTOR'("01000000");
				HEX1 <= STD_LOGIC_VECTOR'("10000010");
			ELSIF P1 = 61 THEN
				HEX0 <= STD_LOGIC_VECTOR'("01111001");
				HEX1 <= STD_LOGIC_VECTOR'("10000010");
			ELSIF P1 = 62 THEN
				HEX0 <= STD_LOGIC_VECTOR'("00100100");
				HEX1 <= STD_LOGIC_VECTOR'("10000010");
			ELSIF P1 = 63 THEN
				HEX0 <= STD_LOGIC_VECTOR'("00110000");
				HEX1 <= STD_LOGIC_VECTOR'("10000010");
			ELSIF P1 = 64 THEN
				HEX0 <= STD_LOGIC_VECTOR'("00011001");
				HEX1 <= STD_LOGIC_VECTOR'("10000010");
			ELSIF P1 = 65 THEN
				HEX0 <= STD_LOGIC_VECTOR'("00010010");
				HEX1 <= STD_LOGIC_VECTOR'("10000010");
			ELSIF P1 = 66 THEN
				HEX0 <= STD_LOGIC_VECTOR'("00000010");
				HEX1 <= STD_LOGIC_VECTOR'("10000010");
			ELSIF P1 = 67 THEN
				HEX0 <= STD_LOGIC_VECTOR'("01111000");
				HEX1 <= STD_LOGIC_VECTOR'("10000010");
			ELSIF P1 = 68 THEN
				HEX0 <= STD_LOGIC_VECTOR'("00000000");
				HEX1 <= STD_LOGIC_VECTOR'("10000010");
			ELSIF P1 = 69 THEN
				HEX0 <= STD_LOGIC_VECTOR'("00011000");
				HEX1 <= STD_LOGIC_VECTOR'("10000010");
			ELSIF P1 = 70 THEN
				HEX0 <= STD_LOGIC_VECTOR'("01000000");
				HEX1 <= STD_LOGIC_VECTOR'("11111000");
			ELSIF P1 = 71 THEN
				HEX0 <= STD_LOGIC_VECTOR'("01111001");
				HEX1 <= STD_LOGIC_VECTOR'("11111000");
			ELSIF P1 = 72 THEN
				HEX0 <= STD_LOGIC_VECTOR'("00100100");
				HEX1 <= STD_LOGIC_VECTOR'("11111000");
			ELSIF P1 = 73 THEN
				HEX0 <= STD_LOGIC_VECTOR'("00110000");
				HEX1 <= STD_LOGIC_VECTOR'("11111000");
			ELSIF P1 = 74 THEN
				HEX0 <= STD_LOGIC_VECTOR'("00011001");
				HEX1 <= STD_LOGIC_VECTOR'("11111000");
			ELSIF P1 = 75 THEN
				HEX0 <= STD_LOGIC_VECTOR'("00010010");
				HEX1 <= STD_LOGIC_VECTOR'("11111000");
			ELSIF P1 = 76 THEN
				HEX0 <= STD_LOGIC_VECTOR'("00000010");
				HEX1 <= STD_LOGIC_VECTOR'("11111000");
			ELSIF P1 = 77 THEN
				HEX0 <= STD_LOGIC_VECTOR'("01111000");
				HEX1 <= STD_LOGIC_VECTOR'("11111000");
			ELSIF P1 = 78 THEN
				HEX0 <= STD_LOGIC_VECTOR'("00000000");
				HEX1 <= STD_LOGIC_VECTOR'("11111000");
			ELSIF P1 = 79 THEN
				HEX0 <= STD_LOGIC_VECTOR'("00011000");
				HEX1 <= STD_LOGIC_VECTOR'("11111000");
			ELSIF P1 = 80 THEN
				HEX0 <= STD_LOGIC_VECTOR'("01000000");
				HEX1 <= STD_LOGIC_VECTOR'("10000000");
			ELSIF P1 = 81 THEN
				HEX0 <= STD_LOGIC_VECTOR'("01111001");
				HEX1 <= STD_LOGIC_VECTOR'("10000000");
			ELSIF P1 = 82 THEN
				HEX0 <= STD_LOGIC_VECTOR'("00100100");
				HEX1 <= STD_LOGIC_VECTOR'("10000000");
			ELSIF P1 = 83 THEN
				HEX0 <= STD_LOGIC_VECTOR'("00110000");
				HEX1 <= STD_LOGIC_VECTOR'("10000000");
			ELSIF P1 = 84 THEN
				HEX0 <= STD_LOGIC_VECTOR'("00011001");
				HEX1 <= STD_LOGIC_VECTOR'("10000000");
			ELSIF P1 = 85 THEN
				HEX0 <= STD_LOGIC_VECTOR'("00010010");
				HEX1 <= STD_LOGIC_VECTOR'("10000000");
			ELSIF P1 = 86 THEN
				HEX0 <= STD_LOGIC_VECTOR'("00000010");
				HEX1 <= STD_LOGIC_VECTOR'("10000000");
			ELSIF P1 = 87 THEN
				HEX0 <= STD_LOGIC_VECTOR'("01111000");
				HEX1 <= STD_LOGIC_VECTOR'("10000000");
			ELSIF P1 = 88 THEN
				HEX0 <= STD_LOGIC_VECTOR'("00000000");
				HEX1 <= STD_LOGIC_VECTOR'("10000000");
			ELSIF P1 = 89 THEN
				HEX0 <= STD_LOGIC_VECTOR'("00011000");
				HEX1 <= STD_LOGIC_VECTOR'("10000000");
			ELSIF P1 = 90 THEN
				HEX0 <= STD_LOGIC_VECTOR'("01000000");
				HEX1 <= STD_LOGIC_VECTOR'("10011000");
			ELSIF P1 = 91 THEN
				HEX0 <= STD_LOGIC_VECTOR'("01111001");
				HEX1 <= STD_LOGIC_VECTOR'("10011000");
			ELSIF P1 = 92 THEN
				HEX0 <= STD_LOGIC_VECTOR'("00100100");
				HEX1 <= STD_LOGIC_VECTOR'("10011000");
			ELSIF P1 = 93 THEN
				HEX0 <= STD_LOGIC_VECTOR'("00110000");
				HEX1 <= STD_LOGIC_VECTOR'("10011000");
			ELSIF P1 = 94 THEN
				HEX0 <= STD_LOGIC_VECTOR'("00011001");
				HEX1 <= STD_LOGIC_VECTOR'("10011000");
			ELSIF P1 = 95 THEN
				HEX0 <= STD_LOGIC_VECTOR'("00010010");
				HEX1 <= STD_LOGIC_VECTOR'("10011000");
			ELSIF P1 = 96 THEN
				HEX0 <= STD_LOGIC_VECTOR'("00000010");
				HEX1 <= STD_LOGIC_VECTOR'("10011000");
			ELSIF P1 = 97 THEN
				HEX0 <= STD_LOGIC_VECTOR'("01111000");
				HEX1 <= STD_LOGIC_VECTOR'("10011000");
			ELSIF P1 = 98 THEN
				HEX0 <= STD_LOGIC_VECTOR'("00000000");
				HEX1 <= STD_LOGIC_VECTOR'("10011000");
			ELSIF P1 = 99 THEN
				HEX0 <= STD_LOGIC_VECTOR'("00011000");
				HEX1 <= STD_LOGIC_VECTOR'("10011000");
			ELSE
				HEX0 <= STD_LOGIC_VECTOR'("11111111");
				HEX1 <= STD_LOGIC_VECTOR'("11111111");
			END IF;
			
		END IF;
			
		IF K <= '1' AND L <= '0' THEN
			IF RSEST = '1' THEN
				IF FALLING_EDGE(MIC_SEC_FLIP) THEN
					P2 := P2 + 1;
				END IF;
			ELSE
				P2 := 0;
			END IF;
		ELSIF K <= '0' AND L <= '1' THEN
			IF RSEST = '1' THEN
					P2 := P2;
			ELSE
				P2 := 0;
			END IF;
		END IF;
		
		IF (P2 = 60) THEN
			SEC_FLIP <= '0';
			P2 :=   0;
		ELSE
			SEC_FLIP <= '1';
			P2 :=   P2;
		END IF;
		
		IF    P2 = 0 THEN
			HEX2 <= STD_LOGIC_VECTOR'("01000000");
			HEX3 <= STD_LOGIC_VECTOR'("11000000");
		ELSIF P2 = 1 THEN
			HEX2 <= STD_LOGIC_VECTOR'("01111001");
			HEX3 <= STD_LOGIC_VECTOR'("11000000");
		ELSIF P2 = 2 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00100100");
			HEX3 <= STD_LOGIC_VECTOR'("11000000");
		ELSIF P2 = 3 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00110000");
			HEX3 <= STD_LOGIC_VECTOR'("11000000");
		ELSIF P2 = 4 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00011001");
			HEX3 <= STD_LOGIC_VECTOR'("11000000");
		ELSIF P2 = 5 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00010010");
			HEX3 <= STD_LOGIC_VECTOR'("11000000");
		ELSIF P2 = 6 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00000010");
			HEX3 <= STD_LOGIC_VECTOR'("11000000");
		ELSIF P2 = 7 THEN
			HEX2 <= STD_LOGIC_VECTOR'("01111000");
			HEX3 <= STD_LOGIC_VECTOR'("11000000");
		ELSIF P2 = 8 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00000000");
			HEX3 <= STD_LOGIC_VECTOR'("11000000");
		ELSIF P2 = 9 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00011000");
			HEX3 <= STD_LOGIC_VECTOR'("11000000");
		ELSIF P2 = 10 THEN
			HEX2 <= STD_LOGIC_VECTOR'("01000000");
			HEX3 <= STD_LOGIC_VECTOR'("11111001");
		ELSIF P2 = 11 THEN
			HEX2 <= STD_LOGIC_VECTOR'("01111001");
			HEX3 <= STD_LOGIC_VECTOR'("11111001");
		ELSIF P2 = 12 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00100100");
			HEX3 <= STD_LOGIC_VECTOR'("11111001");
		ELSIF P2 = 13 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00110000");
			HEX3 <= STD_LOGIC_VECTOR'("11111001");
		ELSIF P2 = 14 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00011001");
			HEX3 <= STD_LOGIC_VECTOR'("11111001");
		ELSIF P2 = 15 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00010010");
			HEX3 <= STD_LOGIC_VECTOR'("11111001");
		ELSIF P2 = 16 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00000010");
			HEX3 <= STD_LOGIC_VECTOR'("11111001");
		ELSIF P2 = 17 THEN
			HEX2 <= STD_LOGIC_VECTOR'("01111000");
			HEX3 <= STD_LOGIC_VECTOR'("11111001");
		ELSIF P2 = 18 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00000000");
			HEX3 <= STD_LOGIC_VECTOR'("11111001");
		ELSIF P2 = 19 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00011000");
			HEX3 <= STD_LOGIC_VECTOR'("11111001");
		ELSIF P2 = 20 THEN
			HEX2 <= STD_LOGIC_VECTOR'("01000000");
			HEX3 <= STD_LOGIC_VECTOR'("10100100");
		ELSIF P2 = 21 THEN
			HEX2 <= STD_LOGIC_VECTOR'("01111001");
			HEX3 <= STD_LOGIC_VECTOR'("10100100");
		ELSIF P2 = 22 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00100100");
			HEX3 <= STD_LOGIC_VECTOR'("10100100");
		ELSIF P2 = 23 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00110000");
			HEX3 <= STD_LOGIC_VECTOR'("10100100");
		ELSIF P2 = 24 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00011001");
			HEX3 <= STD_LOGIC_VECTOR'("10100100");
		ELSIF P2 = 25 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00010010");
			HEX3 <= STD_LOGIC_VECTOR'("10100100");
		ELSIF P2 = 26 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00000010");
			HEX3 <= STD_LOGIC_VECTOR'("10100100");
		ELSIF P2 = 27 THEN
			HEX2 <= STD_LOGIC_VECTOR'("01111000");
			HEX3 <= STD_LOGIC_VECTOR'("10100100");
		ELSIF P2 = 28 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00000000");
			HEX3 <= STD_LOGIC_VECTOR'("10100100");
		ELSIF P2 = 29 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00011000");
			HEX3 <= STD_LOGIC_VECTOR'("10100100");
		ELSIF P2 = 30 THEN
			HEX2 <= STD_LOGIC_VECTOR'("01000000");
			HEX3 <= STD_LOGIC_VECTOR'("10110000");
		ELSIF P2 = 31 THEN
			HEX2 <= STD_LOGIC_VECTOR'("01111001");
			HEX3 <= STD_LOGIC_VECTOR'("10110000");
		ELSIF P2 = 32 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00100100");
			HEX3 <= STD_LOGIC_VECTOR'("10110000");
		ELSIF P2 = 33 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00110000");
			HEX3 <= STD_LOGIC_VECTOR'("10110000");
		ELSIF P2 = 34 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00011001");
			HEX3 <= STD_LOGIC_VECTOR'("10110000");
		ELSIF P2 = 35 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00010010");
			HEX3 <= STD_LOGIC_VECTOR'("10110000");
		ELSIF P2 = 36 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00000010");
			HEX3 <= STD_LOGIC_VECTOR'("10110000");
		ELSIF P2 = 37 THEN
			HEX2 <= STD_LOGIC_VECTOR'("01111000");
			HEX3 <= STD_LOGIC_VECTOR'("10110000");
		ELSIF P2 = 38 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00000000");
			HEX3 <= STD_LOGIC_VECTOR'("10110000");
		ELSIF P2 = 39 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00011000");
			HEX3 <= STD_LOGIC_VECTOR'("10110000");
		ELSIF P2 = 40 THEN
			HEX2 <= STD_LOGIC_VECTOR'("01000000");
			HEX3 <= STD_LOGIC_VECTOR'("10011001");
		ELSIF P2 = 41 THEN
			HEX2 <= STD_LOGIC_VECTOR'("01111001");
			HEX3 <= STD_LOGIC_VECTOR'("10011001");
		ELSIF P2 = 42 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00100100");
			HEX3 <= STD_LOGIC_VECTOR'("10011001");
		ELSIF P2 = 43 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00110000");
			HEX3 <= STD_LOGIC_VECTOR'("10011001");
		ELSIF P2 = 44 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00011001");
			HEX3 <= STD_LOGIC_VECTOR'("10011001");
		ELSIF P2 = 45 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00010010");
			HEX3 <= STD_LOGIC_VECTOR'("10011001");
		ELSIF P2 = 46 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00000010");
			HEX3 <= STD_LOGIC_VECTOR'("10011001");
		ELSIF P2 = 47 THEN
			HEX2 <= STD_LOGIC_VECTOR'("01111000");
			HEX3 <= STD_LOGIC_VECTOR'("10011001");
		ELSIF P2 = 48 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00000000");
			HEX3 <= STD_LOGIC_VECTOR'("10011001");
		ELSIF P2 = 49 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00011000");
			HEX3 <= STD_LOGIC_VECTOR'("10011001");
		ELSIF P2 = 50 THEN
			HEX2 <= STD_LOGIC_VECTOR'("01000000");
			HEX3 <= STD_LOGIC_VECTOR'("10010010");
		ELSIF P2 = 51 THEN
			HEX2 <= STD_LOGIC_VECTOR'("01111001");
			HEX3 <= STD_LOGIC_VECTOR'("10010010");
		ELSIF P2 = 52 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00100100");
			HEX3 <= STD_LOGIC_VECTOR'("10010010");
		ELSIF P2 = 53 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00110000");
			HEX3 <= STD_LOGIC_VECTOR'("10010010");
		ELSIF P2 = 54 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00011001");
			HEX3 <= STD_LOGIC_VECTOR'("10010010");
		ELSIF P2 = 55 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00010010");
			HEX3 <= STD_LOGIC_VECTOR'("10010010");
		ELSIF P2 = 56 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00000010");
			HEX3 <= STD_LOGIC_VECTOR'("10010010");
		ELSIF P2 = 57 THEN
			HEX2 <= STD_LOGIC_VECTOR'("01111000");
			HEX3 <= STD_LOGIC_VECTOR'("10010010");
		ELSIF P2 = 58 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00000000");
			HEX3 <= STD_LOGIC_VECTOR'("10010010");
		ELSIF P2 = 59 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00011000");
			HEX3 <= STD_LOGIC_VECTOR'("10010010");
		ELSE
			HEX2 <= STD_LOGIC_VECTOR'("11111111");
			HEX3 <= STD_LOGIC_VECTOR'("11111111");
		END IF;
		
		IF K <= '1' AND L <= '0' THEN
			IF RSEST = '1' THEN
				IF FALLING_EDGE(SEC_FLIP) THEN
					P3 := P3 + 1;
				END IF;
			ELSE
				P3 := 0;
			END IF;
		ELSIF K <= '0' AND L <= '1' THEN
			IF RSEST = '1' THEN
				P3 := P3;
			ELSE
				P3 := 0;
			END IF;
		END IF;
		
		IF (P3 = 60) THEN
			P3 := 0;
		ELSE
			P3 := P3;
		END IF;
		
		IF    P3 = 0 THEN
			HEX4 <= STD_LOGIC_VECTOR'("01000000");
			HEX5 <= STD_LOGIC_VECTOR'("11000000");
		ELSIF P3 = 1 THEN
			HEX4 <= STD_LOGIC_VECTOR'("01111001");
			HEX5 <= STD_LOGIC_VECTOR'("11000000");
		ELSIF P3 = 2 THEN
			HEX4 <= STD_LOGIC_VECTOR'("00100100");
			HEX5 <= STD_LOGIC_VECTOR'("11000000");
		ELSIF P3 = 3 THEN
			HEX4 <= STD_LOGIC_VECTOR'("00110000");
			HEX5 <= STD_LOGIC_VECTOR'("11000000");
		ELSIF P3 = 4 THEN
			HEX4 <= STD_LOGIC_VECTOR'("00011001");
			HEX5 <= STD_LOGIC_VECTOR'("11000000");
		ELSIF P3 = 5 THEN
			HEX4 <= STD_LOGIC_VECTOR'("00010010");
			HEX5 <= STD_LOGIC_VECTOR'("11000000");
		ELSIF P3 = 6 THEN
			HEX4 <= STD_LOGIC_VECTOR'("00000010");
			HEX5 <= STD_LOGIC_VECTOR'("11000000");
		ELSIF P3 = 7 THEN
			HEX4 <= STD_LOGIC_VECTOR'("01111000");
			HEX5 <= STD_LOGIC_VECTOR'("11000000");
		ELSIF P3 = 8 THEN
			HEX4 <= STD_LOGIC_VECTOR'("00000000");
			HEX5 <= STD_LOGIC_VECTOR'("11000000");
		ELSIF P3 = 9 THEN
			HEX4 <= STD_LOGIC_VECTOR'("00011000");
			HEX5 <= STD_LOGIC_VECTOR'("11000000");
		ELSIF P3 = 10 THEN
			HEX4 <= STD_LOGIC_VECTOR'("01000000");
			HEX5 <= STD_LOGIC_VECTOR'("11111001");
		ELSIF P3 = 11 THEN
			HEX4 <= STD_LOGIC_VECTOR'("01111001");
			HEX5 <= STD_LOGIC_VECTOR'("11111001");
		ELSIF P3 = 12 THEN
			HEX4 <= STD_LOGIC_VECTOR'("00100100");
			HEX5 <= STD_LOGIC_VECTOR'("11111001");
		ELSIF P3 = 13 THEN
			HEX4 <= STD_LOGIC_VECTOR'("00110000");
			HEX5 <= STD_LOGIC_VECTOR'("11111001");
		ELSIF P3 = 14 THEN
			HEX4 <= STD_LOGIC_VECTOR'("00011001");
			HEX5 <= STD_LOGIC_VECTOR'("11111001");
		ELSIF P3 = 15 THEN
			HEX4 <= STD_LOGIC_VECTOR'("00010010");
			HEX5 <= STD_LOGIC_VECTOR'("11111001");
		ELSIF P3 = 16 THEN
			HEX4 <= STD_LOGIC_VECTOR'("00000010");
			HEX5 <= STD_LOGIC_VECTOR'("11111001");
		ELSIF P3 = 17 THEN
			HEX4 <= STD_LOGIC_VECTOR'("01111000");
			HEX5 <= STD_LOGIC_VECTOR'("11111001");
		ELSIF P3 = 18 THEN
			HEX4 <= STD_LOGIC_VECTOR'("00000000");
			HEX5 <= STD_LOGIC_VECTOR'("11111001");
		ELSIF P3 = 19 THEN
			HEX4 <= STD_LOGIC_VECTOR'("00011000");
			HEX5 <= STD_LOGIC_VECTOR'("11111001");
		ELSIF P3 = 20 THEN
			HEX4 <= STD_LOGIC_VECTOR'("01000000");
			HEX5 <= STD_LOGIC_VECTOR'("10100100");
		ELSIF P3 = 21 THEN
			HEX4 <= STD_LOGIC_VECTOR'("01111001");
			HEX5 <= STD_LOGIC_VECTOR'("10100100");
		ELSIF P3 = 22 THEN
			HEX4 <= STD_LOGIC_VECTOR'("00100100");
			HEX5 <= STD_LOGIC_VECTOR'("10100100");
		ELSIF P3 = 23 THEN
			HEX4 <= STD_LOGIC_VECTOR'("00110000");
			HEX5 <= STD_LOGIC_VECTOR'("10100100");
		ELSIF P3 = 24 THEN
			HEX4 <= STD_LOGIC_VECTOR'("00011001");
			HEX5 <= STD_LOGIC_VECTOR'("10100100");
		ELSIF P3 = 25 THEN
			HEX4 <= STD_LOGIC_VECTOR'("00010010");
			HEX5 <= STD_LOGIC_VECTOR'("10100100");
		ELSIF P3 = 26 THEN
			HEX4 <= STD_LOGIC_VECTOR'("00000010");
			HEX5 <= STD_LOGIC_VECTOR'("10100100");
		ELSIF P3 = 27 THEN
			HEX4 <= STD_LOGIC_VECTOR'("01111000");
			HEX5 <= STD_LOGIC_VECTOR'("10100100");
		ELSIF P3 = 28 THEN
			HEX4 <= STD_LOGIC_VECTOR'("00000000");
			HEX5 <= STD_LOGIC_VECTOR'("10100100");
		ELSIF P3 = 29 THEN
			HEX4 <= STD_LOGIC_VECTOR'("00011000");
			HEX5 <= STD_LOGIC_VECTOR'("10100100");
		ELSIF P3 = 30 THEN
			HEX4 <= STD_LOGIC_VECTOR'("01000000");
			HEX5 <= STD_LOGIC_VECTOR'("10110000");
		ELSIF P3 = 31 THEN
			HEX4 <= STD_LOGIC_VECTOR'("01111001");
			HEX5 <= STD_LOGIC_VECTOR'("10110000");
		ELSIF P3 = 32 THEN
			HEX4 <= STD_LOGIC_VECTOR'("00100100");
			HEX5 <= STD_LOGIC_VECTOR'("10110000");
		ELSIF P3 = 33 THEN
			HEX4 <= STD_LOGIC_VECTOR'("00110000");
			HEX5 <= STD_LOGIC_VECTOR'("10110000");
		ELSIF P3 = 34 THEN
			HEX4 <= STD_LOGIC_VECTOR'("00011001");
			HEX5 <= STD_LOGIC_VECTOR'("10110000");
		ELSIF P3 = 35 THEN
			HEX4 <= STD_LOGIC_VECTOR'("00010010");
			HEX5 <= STD_LOGIC_VECTOR'("10110000");
		ELSIF P3 = 36 THEN
			HEX4 <= STD_LOGIC_VECTOR'("00000010");
			HEX5 <= STD_LOGIC_VECTOR'("10110000");
		ELSIF P3 = 37 THEN
			HEX4 <= STD_LOGIC_VECTOR'("01111000");
			HEX5 <= STD_LOGIC_VECTOR'("10110000");
		ELSIF P3 = 38 THEN
			HEX4 <= STD_LOGIC_VECTOR'("00000000");
			HEX5 <= STD_LOGIC_VECTOR'("10110000");
		ELSIF P3 = 39 THEN
			HEX4 <= STD_LOGIC_VECTOR'("00011000");
			HEX5 <= STD_LOGIC_VECTOR'("10110000");
		ELSIF P3 = 40 THEN
			HEX4 <= STD_LOGIC_VECTOR'("01000000");
			HEX5 <= STD_LOGIC_VECTOR'("10011001");
		ELSIF P3 = 41 THEN
			HEX4 <= STD_LOGIC_VECTOR'("01111001");
			HEX5 <= STD_LOGIC_VECTOR'("10011001");
		ELSIF P3 = 42 THEN
			HEX4 <= STD_LOGIC_VECTOR'("00100100");
			HEX5 <= STD_LOGIC_VECTOR'("10011001");
		ELSIF P3 = 43 THEN
			HEX4 <= STD_LOGIC_VECTOR'("00110000");
			HEX5 <= STD_LOGIC_VECTOR'("10011001");
		ELSIF P3 = 44 THEN
			HEX4 <= STD_LOGIC_VECTOR'("00011001");
			HEX5 <= STD_LOGIC_VECTOR'("10011001");
		ELSIF P3 = 45 THEN
			HEX4 <= STD_LOGIC_VECTOR'("00010010");
			HEX5 <= STD_LOGIC_VECTOR'("10011001");
		ELSIF P3 = 46 THEN
			HEX4 <= STD_LOGIC_VECTOR'("00000010");
			HEX5 <= STD_LOGIC_VECTOR'("10011001");
		ELSIF P3 = 47 THEN
			HEX4 <= STD_LOGIC_VECTOR'("01111000");
			HEX5 <= STD_LOGIC_VECTOR'("10011001");
		ELSIF P3 = 48 THEN
			HEX4 <= STD_LOGIC_VECTOR'("00000000");
			HEX5 <= STD_LOGIC_VECTOR'("10011001");
		ELSIF P3 = 49 THEN
			HEX4 <= STD_LOGIC_VECTOR'("00011000");
			HEX5 <= STD_LOGIC_VECTOR'("10011001");
		ELSIF P3 = 50 THEN
			HEX4 <= STD_LOGIC_VECTOR'("01000000");
			HEX5 <= STD_LOGIC_VECTOR'("10010010");
		ELSIF P3 = 51 THEN
			HEX4 <= STD_LOGIC_VECTOR'("01111001");
			HEX5 <= STD_LOGIC_VECTOR'("10010010");
		ELSIF P3 = 52 THEN
			HEX4 <= STD_LOGIC_VECTOR'("00100100");
			HEX5 <= STD_LOGIC_VECTOR'("10010010");
		ELSIF P3 = 53 THEN
			HEX4 <= STD_LOGIC_VECTOR'("00110000");
			HEX5 <= STD_LOGIC_VECTOR'("10010010");
		ELSIF P3 = 54 THEN
			HEX4 <= STD_LOGIC_VECTOR'("00011001");
			HEX5 <= STD_LOGIC_VECTOR'("10010010");
		ELSIF P3 = 55 THEN
			HEX4 <= STD_LOGIC_VECTOR'("00010010");
			HEX5 <= STD_LOGIC_VECTOR'("10010010");
		ELSIF P3 = 56 THEN
			HEX4 <= STD_LOGIC_VECTOR'("00000010");
			HEX5 <= STD_LOGIC_VECTOR'("10010010");
		ELSIF P3 = 57 THEN
			HEX4 <= STD_LOGIC_VECTOR'("01111000");
			HEX5 <= STD_LOGIC_VECTOR'("10010010");
		ELSIF P3 = 58 THEN
			HEX4 <= STD_LOGIC_VECTOR'("00000000");
			HEX5 <= STD_LOGIC_VECTOR'("10010010");
		ELSIF P3 = 59 THEN
			HEX4 <= STD_LOGIC_VECTOR'("00011000");
			HEX5 <= STD_LOGIC_VECTOR'("10010010");
		ELSE
			HEX4 <= STD_LOGIC_VECTOR'("11111111");
			HEX5 <= STD_LOGIC_VECTOR'("11111111");
		END IF;
		
	END IF;
	
END PROCESS;
END behaviour;